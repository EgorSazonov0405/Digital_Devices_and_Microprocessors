module module_3_lab_2 (
    input logic [3:0] din,
    output logic [3:0] dout
);
// Преобразование из двоичного кода в код Грея выполняется по простому правилу:
//Старший бит кода Грея равен старшему биту двоичного кода
// Каждый следующий бит кода Грея получается как XOR (исключающее ИЛИ) между соответствующим и старшим соседним битом двоичного кода
//
//Преобразование по правилам кода Грея
//
assign dout[3] = din[3];
assign dout[2] = din[3] ^ din[2]; // XOR между битами
assign dout[1] = din[2] ^ din[1];
assign dout[0] = din[1] ^ din[0];

endmodule