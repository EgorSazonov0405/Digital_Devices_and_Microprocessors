module tb_lab92();

logic clk;
logic [7:0] x1;
logic [7:0] x2;
logic [7:0] dout;

lab92 dut (
    .clk(clk),
    .x1(x1),
    .x2(x2),
    .dout(dout)
);
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Test cases
    initial begin
        // Тест 1: Оба положительные, простой случай
        x1 = 8'b0001_0000; // 1.0 в (1,8,4): 16/16 = 1.0
        x2 = 8'b0001_0000; // 1.0 в (1,8,4): 16/16 = 1.0
        #10;
        // Тест 2: Оба положительные, дробные числа
        x1 = 8'b0000_1000; // 0.5 в (1,8,4): 8/16 = 0.5
        x2 = 8'b0000_1000; // 0.5 в (1,8,4): 8/16 = 0.5
        #10;
        // Тест 3: Отрицательное × положительное
        x1 = 8'b1111_0000; // -1.0 в (1,8,4): -16/16 = -1.0
        x2 = 8'b0001_0000; // 1.0 в (1,8,4): 16/16 = 1.0
        #10;
        // Тест 4: Оба отрицательные
        x1 = 8'b1111_0000; // -1.0 в (1,8,4): -16/16 = -1.0
        x2 = 8'b1111_0000; // -1.0 в (1,8,4): -16/16 = -1.0
        #10;
        // Тест 5: Максимальные положительные значения
        x1 = 8'b0111_1111; // 7.9375 в (1,8,4): 127/16 ≈ 7.9375
        x2 = 8'b0000_0001; // 0.0625 в (1,8,4): 1/16 = 0.0625
        #10;        
        // Тест 6: Переполнение (без насыщения)
        x1 = 8'b0111_0000; // 7.0 в (1,8,4): 112/16 = 7.0
        x2 = 8'b0111_0000; // 7.0 в (1,8,4): 112/16 = 7.0
        #10;
        // Тест 7: Нулевые значения
        x1 = 8'b0000_0000; // 0.0
        x2 = 8'b0000_0000; // 0.0
        #10;
        $finish;
    end
endmodule