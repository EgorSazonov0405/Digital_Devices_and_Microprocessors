module module_2_lab_2 (
    input logic [7:0] din,
    output logic [3:0] dout
);
assign dout = (din == 8'b00000001) ? 4'b0000: // только 0
              (din == 8'b00000010) ? 4'b0001: // только 1
              (din == 8'b00000100) ? 4'b0010: // только 2
              (din == 8'b00001000) ? 4'b0011: // только 3
              (din == 8'b00010000) ? 4'b0100: // только 4                                    
              (din == 8'b00100000) ? 4'b0101: // только 5
              (din == 8'b01000000) ? 4'b0110: // только 6
              (din == 8'b1000000) ? 4'b0111: // только 7
              4'b1000; // все остальные случаи - ошибка!                           
//
// ВТОРОЙ ВАРИАНТ РЕШЕНИЯ
//
// always_comb begin
//     case (din)
//         8'b00000001: dout = 4'b0000;
//         8'b00000010: dout = 4'b0001;
//         8'b00000100: dout = 4'b0010;
//         8'b00001000: dout = 4'b0011;
//         8'b00010000: dout = 4'b0100;
//         8'b00100000: dout = 4'b0101;
//         8'b01000000: dout = 4'b0110;
//         8'b10000000: dout = 4'b0111;
//         default:     dout = 4'b1000; // Обработка всех остальных случаев
//     endcase
// end

endmodule