module tb_lab91();

logic clk;
logic [15:0] x1;
logic [7:0] x2;
logic [20:0] dout;

// Instantiate DUT
lab91 dut (
    .clk(clk),
    .x1(x1),
    .x2(x2),
    .dout(dout)
);
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Tests
    initial begin    
        // Тест 1: Оба положительные
        x1 = 16'b0000_0000_1000_0000; // 0.5 в (1,16,8): 128/256 = 0.5
        x2 = 8'b0000_1000;           // 0.03125 в (1,8,12): 8/4096 = 0.001953125
        #10;
        // Тест 2: Оба отрицательные
        x1 = 16'b1111_1111_1000_0000; // -0.5 в (1,16,8): -128/256 = -0.5
        x2 = 8'b1111_1000;           // -0.03125 в (1,8,12): -8/4096 = -0.001953125
        #10;
        // Тест 3: Разные знаки (x1 положительный, x2 отрицательный)
        x1 = 16'b0000_0000_1100_0000; // 0.75 в (1,16,8): 192/256 = 0.75
        x2 = 8'b1111_0000;           // -0.0625 в (1,8,12): -16/4096 = -0.00390625
        #10;
        // Тест 4: Разные знаки (x1 отрицательный, x2 положительный)
        x1 = 16'b1111_1111_0100_0000; // -0.75 в (1,16,8): -192/256 = -0.75
        x2 = 8'b0001_0000;           // 0.0625 в (1,8,12): 16/4096 = 0.00390625
        #10;
        // Тест 5: Граничные значения
        x1 = 16'b0111_1111_1111_1111; // Максимальное положительное: 32767/256 ≈ 127.996
        x2 = 8'b0111_1111;           // Максимальное положительное: 127/4096 ≈ 0.031
        #10;
        // Тест 6: Нулевые значения
        x1 = 16'b0000_0000_0000_0000; // 0
        x2 = 8'b0000_0000;           // 0
        #10;
        $finish;
    end
endmodule