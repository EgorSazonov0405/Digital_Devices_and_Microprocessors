module module_4_lab_2 (
    input logic [4 : 0] din, // 5 разряд. двоичный код
    output logic [6 : 0] dout, // 7-сегментный код
    output logic [3 : 0] an // Управление анодами
);
// Приоритетный шифратор — это цифровая схема, которая определяет позицию старшего (наивысшего) установленного бита во входном слове.

// Активация только правого индикатора
assign an = 4'b1110;

assign dout = (din[4] == 1'b1) ? ~7'b1100110 : // 4 - log2 от чисел диапазона [16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31] 
              (din[3] == 1'b1) ? ~7'b1001111 : // 3 - log2 от чисел диапазона [8, 9, 10, 11, 12, 13, 14, 15] 
              (din[2] == 1'b1) ? ~7'b1011011 : // 2 - log2 от чисел диапазона [4, 5, 6, 7] 
              (din[1] == 1'b1) ? ~7'b0000110 : // 1 - log2 от чисел диапазона [2, 3]
              (din[0] == 1'b1) ? ~7'b0111111 : // 0 - log2(1)
              ~7'b0111111                      // 0 - log2(0)

endmodule