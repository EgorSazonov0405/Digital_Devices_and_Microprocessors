module module_4_lab_2 (
    input logic [3 : 0] din, // 4 разряд. двоичный код
    output logic [6 : 0] dout, // 7-сегментный код
    output logic [3 : 0] an // Управление анодами
);
// Активация только правого индикатора
assign an = 4'b1110;
// Преобразование двоичного кода в 7-сегментный с инверсией
assign dout = (din == 4'b0000) ? ~7'b0111111 : // 0
              (din == 4'b0001) ? ~7'b0000110 : // 1
              (din == 4'b0010) ? ~7'b1011011 : // 2
              (din == 4'b0011) ? ~7'b1001111 : // 3
              (din == 4'b0100) ? ~7'b1100110 : // 4
              (din == 4'b0101) ? ~7'b1101101 : // 5
              (din == 4'b0110) ? ~7'b1111101 : // 6
              (din == 4'b0111) ? ~7'b0000111 : // 7
              (din == 4'b1000) ? ~7'b1111111 : // 8
              (din == 4'b1001) ? ~7'b1101111 : // 9
              (din == 4'b1010) ? ~7'b1110111 : // 10 - A
              (din == 4'b1011) ? ~7'b1111100 : // 11 - B
              (din == 4'b1100) ? ~7'b0111001 : // 12 - C
              (din == 4'b1101) ? ~7'b1011110 : // 13 - D
              (din == 4'b1110) ? ~7'b1111001 : // 14 - E
              ~7'b1110001; // 15 - F

endmodule