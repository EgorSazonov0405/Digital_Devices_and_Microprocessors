// Блок, выполняющий циклический сдвиг четырехразрядного числа влево на два разряда
module lab43 (
    input logic [3 : 0] x,
    output logic [7 : 0] y
);

assign y[3:0] = x;
assign y[7:4] = {x[1:0], x[3:2]}; // сдвиг на 2 элемента влево

endmodule