module tb_lab93();

    logic clk;
    logic [7:0] x1;
    logic [7:0] x2;
    logic [7:0] dout;

    lab93 dut (
        .clk(clk),
        .x1(x1),
        .x2(x2),
        .dout(dout)
    );

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Test cases
    initial begin
        // Тест 1: Простой случай, без насыщения
        x1 = 8'b0001_0000; // +1.0
        x2 = 8'b0001_0000; // +1.0
        #10;
        // Тест 2: Округление в большую сторону
        x1 = 8'b0000_1000; // 0.5
        x2 = 8'b0000_1001; // 0.5625 (9/16)
        #10;
        // Тест 3: Округление в меньшую сторону
        x1 = 8'b0000_1000; // 0.5
        x2 = 8'b0000_0111; // 0.4375 (7/16)
        #10;
        // Тест 4: Положительное насыщение
        x1 = 8'b0111_0000; // 7.0
        x2 = 8'b0111_0000; // 7.0
        #10;
        // Тест 5: Отрицательное насыщение
        x1 = 8'b1001_0000; // -7.0
        x2 = 8'b1001_0000; // -7.0
        #10;
        // Тест 6: Граничный случай - чуть ниже насыщения
        x1 = 8'b0110_0000; // 6.0
        x2 = 8'b0110_0000; // 6.0
        #10;
        // Тест 7: Отрицательное × положительное с насыщением
        x1 = 8'b1000_0000; // -8.0
        x2 = 8'b0111_0000; // 7.0
        #10;  
        // Тест 8: Проверка округления с отрицательными числами
        x1 = 8'b1111_1000; // -0.5
        x2 = 8'b1111_1001; // -0.4375
        #10;
        $finish;
    end
endmodule